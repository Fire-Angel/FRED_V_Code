`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    23:19:23 02/27/2014 
// Design Name: 
// Module Name:    LoadMSK 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module LoadMSK( clk,  MSK, reset, mem_out);
input clk; 
input reset; 
input wire signed [15:0] MSK ;
output wire signed [15:0] mem_out;  
reg signed [15:0] b [0:199];
reg [7:0] i = 0;
reg signed [19:0] temp;
reg signed [29:0] accumulator = 30'b0000000000000000000000000000000;
reg signed [15:0] zero = 16'b0110011100011101;
reg signed [15:0] one  = 16'b0110011100011101;
assign mem_out = accumulator [29:14];

	 always @(posedge clk) begin
	 if (reset == 1'b1) begin 
	 accumulator = 30'b0000000000000000000000000000000;
	 end 
	 else begin 
	    temp = zero * MSK;
		 accumulator = accumulator + temp;
end		 
		 if (i << 199) begin 
      b[i][0] <= MSK[0];
		b[i][1] <= MSK[1];
		b[i][2] <= MSK[2];
		b[i][3] <= MSK[3];
		b[i][4] <= MSK[4];
		b[i][5] <= MSK[5];
		b[i][6] <= MSK[6];
		b[i][7] <= MSK[7];
		b[i][8] <= MSK[8];
		b[i][9] <= MSK[9];
		b[i][10] <= MSK[10];
		b[i][11] <= MSK[11];
		b[i][12] <= MSK[12];
		b[i][13] <= MSK[13];
		b[i][14] <= MSK[14];
		b[i][15] <= MSK[15];
		end
	
		else if (i == 199) begin 
      b[0][0] <= MSK[0];
		b[0][1] <= MSK[1];
		b[0][2] <= MSK[2];
		b[0][3] <= MSK[3];
		b[0][4] <= MSK[4];
		b[0][5] <= MSK[5];
		b[0][6] <= MSK[6];
		b[0][7] <= MSK[7];
		b[0][8] <= MSK[8];
		b[0][9] <= MSK[9];
		b[0][10] <= MSK[10];
		b[0][11] <= MSK[11];
		b[0][12] <= MSK[12];
		b[0][13] <= MSK[13];
		b[0][14] <= MSK[14];
		b[0][15] <= MSK[15];
{b[1][0], b[1][1],b[1][2],b[1][3],b[1][4],b[1][5],b[1][6],b[1][7],b[1][8],b[1][9],b[1][10],b[1][11],b[1][12],b[1][13],b[1][14],b[1][15]} <= {b[0][0], b[0][1],b[0][2],b[0][3],b[0][4],b[0][5],b[0][6],b[0][7],b[0][8],b[0][9],b[0][10],b[0][11],b[0][12],b[0][13],b[0][14],b[0][15]}; 
{b[2][0], b[2][1],b[2][2],b[2][3],b[2][4],b[2][5],b[2][6],b[2][7],b[2][8],b[2][9],b[2][10],b[2][11],b[2][12],b[2][13],b[2][14],b[2][15]} <= {b[1][0], b[1][1],b[1][2],b[1][3],b[1][4],b[1][5],b[1][6],b[1][7],b[1][8],b[1][9],b[1][10],b[1][11],b[1][12],b[1][13],b[1][14],b[1][15]}; 
{b[3][0], b[3][1],b[3][2],b[3][3],b[3][4],b[3][5],b[3][6],b[3][7],b[3][8],b[3][9],b[3][10],b[3][11],b[3][12],b[3][13],b[3][14],b[3][15]} <= {b[2][0], b[2][1],b[2][2],b[2][3],b[2][4],b[2][5],b[2][6],b[2][7],b[2][8],b[2][9],b[2][10],b[2][11],b[2][12],b[2][13],b[2][14],b[2][15]}; 
{b[4][0], b[4][1],b[4][2],b[4][3],b[4][4],b[4][5],b[4][6],b[4][7],b[4][8],b[4][9],b[4][10],b[4][11],b[4][12],b[4][13],b[4][14],b[4][15]} <= {b[3][0], b[3][1],b[3][2],b[3][3],b[3][4],b[3][5],b[3][6],b[3][7],b[3][8],b[3][9],b[3][10],b[3][11],b[3][12],b[3][13],b[3][14],b[3][15]}; 
{b[5][0], b[5][1],b[5][2],b[5][3],b[5][4],b[5][5],b[5][6],b[5][7],b[5][8],b[5][9],b[5][10],b[5][11],b[5][12],b[5][13],b[5][14],b[5][15]} <= {b[4][0], b[4][1],b[4][2],b[4][3],b[4][4],b[4][5],b[4][6],b[4][7],b[4][8],b[4][9],b[4][10],b[4][11],b[4][12],b[4][13],b[4][14],b[4][15]}; 
{b[6][0], b[6][1],b[6][2],b[6][3],b[6][4],b[6][5],b[6][6],b[6][7],b[6][8],b[6][9],b[6][10],b[6][11],b[6][12],b[6][13],b[6][14],b[6][15]} <= {b[5][0], b[5][1],b[5][2],b[5][3],b[5][4],b[5][5],b[5][6],b[5][7],b[5][8],b[5][9],b[5][10],b[5][11],b[5][12],b[5][13],b[5][14],b[5][15]}; 
{b[7][0], b[7][1],b[7][2],b[7][3],b[7][4],b[7][5],b[7][6],b[7][7],b[7][8],b[7][9],b[7][10],b[7][11],b[7][12],b[7][13],b[7][14],b[7][15]} <= {b[6][0], b[6][1],b[6][2],b[6][3],b[6][4],b[6][5],b[6][6],b[6][7],b[6][8],b[6][9],b[6][10],b[6][11],b[6][12],b[6][13],b[6][14],b[6][15]}; 
{b[8][0], b[8][1],b[8][2],b[8][3],b[8][4],b[8][5],b[8][6],b[8][7],b[8][8],b[8][9],b[8][10],b[8][11],b[8][12],b[8][13],b[8][14],b[8][15]} <= {b[7][0], b[7][1],b[7][2],b[7][3],b[7][4],b[7][5],b[7][6],b[7][7],b[7][8],b[7][9],b[7][10],b[7][11],b[7][12],b[7][13],b[7][14],b[7][15]}; 
{b[9][0], b[9][1],b[9][2],b[9][3],b[9][4],b[9][5],b[9][6],b[9][7],b[9][8],b[9][9],b[9][10],b[9][11],b[9][12],b[9][13],b[9][14],b[9][15]} <= {b[8][0], b[8][1],b[8][2],b[8][3],b[8][4],b[8][5],b[8][6],b[8][7],b[8][8],b[8][9],b[8][10],b[8][11],b[8][12],b[8][13],b[8][14],b[8][15]}; 
{b[10][0], b[10][1],b[10][2],b[10][3],b[10][4],b[10][5],b[10][6],b[10][7],b[10][8],b[10][9],b[10][10],b[10][11],b[10][12],b[10][13],b[10][14],b[10][15]} <= {b[9][0], b[9][1],b[9][2],b[9][3],b[9][4],b[9][5],b[9][6],b[9][7],b[9][8],b[9][9],b[9][10],b[9][11],b[9][12],b[9][13],b[9][14],b[9][15]}; 
{b[11][0], b[11][1],b[11][2],b[11][3],b[11][4],b[11][5],b[11][6],b[11][7],b[11][8],b[11][9],b[11][10],b[11][11],b[11][12],b[11][13],b[11][14],b[11][15]} <= {b[10][0], b[10][1],b[10][2],b[10][3],b[10][4],b[10][5],b[10][6],b[10][7],b[10][8],b[10][9],b[10][10],b[10][11],b[10][12],b[10][13],b[10][14],b[10][15]}; 
{b[12][0], b[12][1],b[12][2],b[12][3],b[12][4],b[12][5],b[12][6],b[12][7],b[12][8],b[12][9],b[12][10],b[12][11],b[12][12],b[12][13],b[12][14],b[12][15]} <= {b[11][0], b[11][1],b[11][2],b[11][3],b[11][4],b[11][5],b[11][6],b[11][7],b[11][8],b[11][9],b[11][10],b[11][11],b[11][12],b[11][13],b[11][14],b[11][15]}; 
{b[13][0], b[13][1],b[13][2],b[13][3],b[13][4],b[13][5],b[13][6],b[13][7],b[13][8],b[13][9],b[13][10],b[13][11],b[13][12],b[13][13],b[13][14],b[13][15]} <= {b[12][0], b[12][1],b[12][2],b[12][3],b[12][4],b[12][5],b[12][6],b[12][7],b[12][8],b[12][9],b[12][10],b[12][11],b[12][12],b[12][13],b[12][14],b[12][15]}; 
{b[14][0], b[14][1],b[14][2],b[14][3],b[14][4],b[14][5],b[14][6],b[14][7],b[14][8],b[14][9],b[14][10],b[14][11],b[14][12],b[14][13],b[14][14],b[14][15]} <= {b[13][0], b[13][1],b[13][2],b[13][3],b[13][4],b[13][5],b[13][6],b[13][7],b[13][8],b[13][9],b[13][10],b[13][11],b[13][12],b[13][13],b[13][14],b[13][15]}; 
{b[15][0], b[15][1],b[15][2],b[15][3],b[15][4],b[15][5],b[15][6],b[15][7],b[15][8],b[15][9],b[15][10],b[15][11],b[15][12],b[15][13],b[15][14],b[15][15]} <= {b[14][0], b[14][1],b[14][2],b[14][3],b[14][4],b[14][5],b[14][6],b[14][7],b[14][8],b[14][9],b[14][10],b[14][11],b[14][12],b[14][13],b[14][14],b[14][15]}; 
{b[16][0], b[16][1],b[16][2],b[16][3],b[16][4],b[16][5],b[16][6],b[16][7],b[16][8],b[16][9],b[16][10],b[16][11],b[16][12],b[16][13],b[16][14],b[16][15]} <= {b[15][0], b[15][1],b[15][2],b[15][3],b[15][4],b[15][5],b[15][6],b[15][7],b[15][8],b[15][9],b[15][10],b[15][11],b[15][12],b[15][13],b[15][14],b[15][15]}; 
{b[17][0], b[17][1],b[17][2],b[17][3],b[17][4],b[17][5],b[17][6],b[17][7],b[17][8],b[17][9],b[17][10],b[17][11],b[17][12],b[17][13],b[17][14],b[17][15]} <= {b[16][0], b[16][1],b[16][2],b[16][3],b[16][4],b[16][5],b[16][6],b[16][7],b[16][8],b[16][9],b[16][10],b[16][11],b[16][12],b[16][13],b[16][14],b[16][15]}; 
{b[18][0], b[18][1],b[18][2],b[18][3],b[18][4],b[18][5],b[18][6],b[18][7],b[18][8],b[18][9],b[18][10],b[18][11],b[18][12],b[18][13],b[18][14],b[18][15]} <= {b[17][0], b[17][1],b[17][2],b[17][3],b[17][4],b[17][5],b[17][6],b[17][7],b[17][8],b[17][9],b[17][10],b[17][11],b[17][12],b[17][13],b[17][14],b[17][15]}; 
{b[19][0], b[19][1],b[19][2],b[19][3],b[19][4],b[19][5],b[19][6],b[19][7],b[19][8],b[19][9],b[19][10],b[19][11],b[19][12],b[19][13],b[19][14],b[19][15]} <= {b[18][0], b[18][1],b[18][2],b[18][3],b[18][4],b[18][5],b[18][6],b[18][7],b[18][8],b[18][9],b[18][10],b[18][11],b[18][12],b[18][13],b[18][14],b[18][15]}; 
{b[20][0], b[20][1],b[20][2],b[20][3],b[20][4],b[20][5],b[20][6],b[20][7],b[20][8],b[20][9],b[20][10],b[20][11],b[20][12],b[20][13],b[20][14],b[20][15]} <= {b[19][0], b[19][1],b[19][2],b[19][3],b[19][4],b[19][5],b[19][6],b[19][7],b[19][8],b[19][9],b[19][10],b[19][11],b[19][12],b[19][13],b[19][14],b[19][15]}; 
{b[21][0], b[21][1],b[21][2],b[21][3],b[21][4],b[21][5],b[21][6],b[21][7],b[21][8],b[21][9],b[21][10],b[21][11],b[21][12],b[21][13],b[21][14],b[21][15]} <= {b[20][0], b[20][1],b[20][2],b[20][3],b[20][4],b[20][5],b[20][6],b[20][7],b[20][8],b[20][9],b[20][10],b[20][11],b[20][12],b[20][13],b[20][14],b[20][15]}; 
{b[22][0], b[22][1],b[22][2],b[22][3],b[22][4],b[22][5],b[22][6],b[22][7],b[22][8],b[22][9],b[22][10],b[22][11],b[22][12],b[22][13],b[22][14],b[22][15]} <= {b[21][0], b[21][1],b[21][2],b[21][3],b[21][4],b[21][5],b[21][6],b[21][7],b[21][8],b[21][9],b[21][10],b[21][11],b[21][12],b[21][13],b[21][14],b[21][15]}; 
{b[23][0], b[23][1],b[23][2],b[23][3],b[23][4],b[23][5],b[23][6],b[23][7],b[23][8],b[23][9],b[23][10],b[23][11],b[23][12],b[23][13],b[23][14],b[23][15]} <= {b[22][0], b[22][1],b[22][2],b[22][3],b[22][4],b[22][5],b[22][6],b[22][7],b[22][8],b[22][9],b[22][10],b[22][11],b[22][12],b[22][13],b[22][14],b[22][15]}; 
{b[24][0], b[24][1],b[24][2],b[24][3],b[24][4],b[24][5],b[24][6],b[24][7],b[24][8],b[24][9],b[24][10],b[24][11],b[24][12],b[24][13],b[24][14],b[24][15]} <= {b[23][0], b[23][1],b[23][2],b[23][3],b[23][4],b[23][5],b[23][6],b[23][7],b[23][8],b[23][9],b[23][10],b[23][11],b[23][12],b[23][13],b[23][14],b[23][15]}; 
{b[25][0], b[25][1],b[25][2],b[25][3],b[25][4],b[25][5],b[25][6],b[25][7],b[25][8],b[25][9],b[25][10],b[25][11],b[25][12],b[25][13],b[25][14],b[25][15]} <= {b[24][0], b[24][1],b[24][2],b[24][3],b[24][4],b[24][5],b[24][6],b[24][7],b[24][8],b[24][9],b[24][10],b[24][11],b[24][12],b[24][13],b[24][14],b[24][15]}; 
{b[26][0], b[26][1],b[26][2],b[26][3],b[26][4],b[26][5],b[26][6],b[26][7],b[26][8],b[26][9],b[26][10],b[26][11],b[26][12],b[26][13],b[26][14],b[26][15]} <= {b[25][0], b[25][1],b[25][2],b[25][3],b[25][4],b[25][5],b[25][6],b[25][7],b[25][8],b[25][9],b[25][10],b[25][11],b[25][12],b[25][13],b[25][14],b[25][15]}; 
{b[27][0], b[27][1],b[27][2],b[27][3],b[27][4],b[27][5],b[27][6],b[27][7],b[27][8],b[27][9],b[27][10],b[27][11],b[27][12],b[27][13],b[27][14],b[27][15]} <= {b[26][0], b[26][1],b[26][2],b[26][3],b[26][4],b[26][5],b[26][6],b[26][7],b[26][8],b[26][9],b[26][10],b[26][11],b[26][12],b[26][13],b[26][14],b[26][15]}; 
{b[28][0], b[28][1],b[28][2],b[28][3],b[28][4],b[28][5],b[28][6],b[28][7],b[28][8],b[28][9],b[28][10],b[28][11],b[28][12],b[28][13],b[28][14],b[28][15]} <= {b[27][0], b[27][1],b[27][2],b[27][3],b[27][4],b[27][5],b[27][6],b[27][7],b[27][8],b[27][9],b[27][10],b[27][11],b[27][12],b[27][13],b[27][14],b[27][15]}; 
{b[29][0], b[29][1],b[29][2],b[29][3],b[29][4],b[29][5],b[29][6],b[29][7],b[29][8],b[29][9],b[29][10],b[29][11],b[29][12],b[29][13],b[29][14],b[29][15]} <= {b[28][0], b[28][1],b[28][2],b[28][3],b[28][4],b[28][5],b[28][6],b[28][7],b[28][8],b[28][9],b[28][10],b[28][11],b[28][12],b[28][13],b[28][14],b[28][15]}; 
{b[30][0], b[30][1],b[30][2],b[30][3],b[30][4],b[30][5],b[30][6],b[30][7],b[30][8],b[30][9],b[30][10],b[30][11],b[30][12],b[30][13],b[30][14],b[30][15]} <= {b[29][0], b[29][1],b[29][2],b[29][3],b[29][4],b[29][5],b[29][6],b[29][7],b[29][8],b[29][9],b[29][10],b[29][11],b[29][12],b[29][13],b[29][14],b[29][15]}; 
{b[31][0], b[31][1],b[31][2],b[31][3],b[31][4],b[31][5],b[31][6],b[31][7],b[31][8],b[31][9],b[31][10],b[31][11],b[31][12],b[31][13],b[31][14],b[31][15]} <= {b[30][0], b[30][1],b[30][2],b[30][3],b[30][4],b[30][5],b[30][6],b[30][7],b[30][8],b[30][9],b[30][10],b[30][11],b[30][12],b[30][13],b[30][14],b[30][15]}; 
{b[32][0], b[32][1],b[32][2],b[32][3],b[32][4],b[32][5],b[32][6],b[32][7],b[32][8],b[32][9],b[32][10],b[32][11],b[32][12],b[32][13],b[32][14],b[32][15]} <= {b[31][0], b[31][1],b[31][2],b[31][3],b[31][4],b[31][5],b[31][6],b[31][7],b[31][8],b[31][9],b[31][10],b[31][11],b[31][12],b[31][13],b[31][14],b[31][15]}; 
{b[33][0], b[33][1],b[33][2],b[33][3],b[33][4],b[33][5],b[33][6],b[33][7],b[33][8],b[33][9],b[33][10],b[33][11],b[33][12],b[33][13],b[33][14],b[33][15]} <= {b[32][0], b[32][1],b[32][2],b[32][3],b[32][4],b[32][5],b[32][6],b[32][7],b[32][8],b[32][9],b[32][10],b[32][11],b[32][12],b[32][13],b[32][14],b[32][15]}; 
{b[34][0], b[34][1],b[34][2],b[34][3],b[34][4],b[34][5],b[34][6],b[34][7],b[34][8],b[34][9],b[34][10],b[34][11],b[34][12],b[34][13],b[34][14],b[34][15]} <= {b[33][0], b[33][1],b[33][2],b[33][3],b[33][4],b[33][5],b[33][6],b[33][7],b[33][8],b[33][9],b[33][10],b[33][11],b[33][12],b[33][13],b[33][14],b[33][15]}; 
{b[35][0], b[35][1],b[35][2],b[35][3],b[35][4],b[35][5],b[35][6],b[35][7],b[35][8],b[35][9],b[35][10],b[35][11],b[35][12],b[35][13],b[35][14],b[35][15]} <= {b[34][0], b[34][1],b[34][2],b[34][3],b[34][4],b[34][5],b[34][6],b[34][7],b[34][8],b[34][9],b[34][10],b[34][11],b[34][12],b[34][13],b[34][14],b[34][15]}; 
{b[36][0], b[36][1],b[36][2],b[36][3],b[36][4],b[36][5],b[36][6],b[36][7],b[36][8],b[36][9],b[36][10],b[36][11],b[36][12],b[36][13],b[36][14],b[36][15]} <= {b[35][0], b[35][1],b[35][2],b[35][3],b[35][4],b[35][5],b[35][6],b[35][7],b[35][8],b[35][9],b[35][10],b[35][11],b[35][12],b[35][13],b[35][14],b[35][15]}; 
{b[37][0], b[37][1],b[37][2],b[37][3],b[37][4],b[37][5],b[37][6],b[37][7],b[37][8],b[37][9],b[37][10],b[37][11],b[37][12],b[37][13],b[37][14],b[37][15]} <= {b[36][0], b[36][1],b[36][2],b[36][3],b[36][4],b[36][5],b[36][6],b[36][7],b[36][8],b[36][9],b[36][10],b[36][11],b[36][12],b[36][13],b[36][14],b[36][15]}; 
{b[38][0], b[38][1],b[38][2],b[38][3],b[38][4],b[38][5],b[38][6],b[38][7],b[38][8],b[38][9],b[38][10],b[38][11],b[38][12],b[38][13],b[38][14],b[38][15]} <= {b[37][0], b[37][1],b[37][2],b[37][3],b[37][4],b[37][5],b[37][6],b[37][7],b[37][8],b[37][9],b[37][10],b[37][11],b[37][12],b[37][13],b[37][14],b[37][15]}; 
{b[39][0], b[39][1],b[39][2],b[39][3],b[39][4],b[39][5],b[39][6],b[39][7],b[39][8],b[39][9],b[39][10],b[39][11],b[39][12],b[39][13],b[39][14],b[39][15]} <= {b[38][0], b[38][1],b[38][2],b[38][3],b[38][4],b[38][5],b[38][6],b[38][7],b[38][8],b[38][9],b[38][10],b[38][11],b[38][12],b[38][13],b[38][14],b[38][15]}; 
{b[40][0], b[40][1],b[40][2],b[40][3],b[40][4],b[40][5],b[40][6],b[40][7],b[40][8],b[40][9],b[40][10],b[40][11],b[40][12],b[40][13],b[40][14],b[40][15]} <= {b[39][0], b[39][1],b[39][2],b[39][3],b[39][4],b[39][5],b[39][6],b[39][7],b[39][8],b[39][9],b[39][10],b[39][11],b[39][12],b[39][13],b[39][14],b[39][15]}; 
{b[41][0], b[41][1],b[41][2],b[41][3],b[41][4],b[41][5],b[41][6],b[41][7],b[41][8],b[41][9],b[41][10],b[41][11],b[41][12],b[41][13],b[41][14],b[41][15]} <= {b[40][0], b[40][1],b[40][2],b[40][3],b[40][4],b[40][5],b[40][6],b[40][7],b[40][8],b[40][9],b[40][10],b[40][11],b[40][12],b[40][13],b[40][14],b[40][15]}; 
{b[42][0], b[42][1],b[42][2],b[42][3],b[42][4],b[42][5],b[42][6],b[42][7],b[42][8],b[42][9],b[42][10],b[42][11],b[42][12],b[42][13],b[42][14],b[42][15]} <= {b[41][0], b[41][1],b[41][2],b[41][3],b[41][4],b[41][5],b[41][6],b[41][7],b[41][8],b[41][9],b[41][10],b[41][11],b[41][12],b[41][13],b[41][14],b[41][15]}; 
{b[43][0], b[43][1],b[43][2],b[43][3],b[43][4],b[43][5],b[43][6],b[43][7],b[43][8],b[43][9],b[43][10],b[43][11],b[43][12],b[43][13],b[43][14],b[43][15]} <= {b[42][0], b[42][1],b[42][2],b[42][3],b[42][4],b[42][5],b[42][6],b[42][7],b[42][8],b[42][9],b[42][10],b[42][11],b[42][12],b[42][13],b[42][14],b[42][15]}; 
{b[44][0], b[44][1],b[44][2],b[44][3],b[44][4],b[44][5],b[44][6],b[44][7],b[44][8],b[44][9],b[44][10],b[44][11],b[44][12],b[44][13],b[44][14],b[44][15]} <= {b[43][0], b[43][1],b[43][2],b[43][3],b[43][4],b[43][5],b[43][6],b[43][7],b[43][8],b[43][9],b[43][10],b[43][11],b[43][12],b[43][13],b[43][14],b[43][15]}; 
{b[45][0], b[45][1],b[45][2],b[45][3],b[45][4],b[45][5],b[45][6],b[45][7],b[45][8],b[45][9],b[45][10],b[45][11],b[45][12],b[45][13],b[45][14],b[45][15]} <= {b[44][0], b[44][1],b[44][2],b[44][3],b[44][4],b[44][5],b[44][6],b[44][7],b[44][8],b[44][9],b[44][10],b[44][11],b[44][12],b[44][13],b[44][14],b[44][15]}; 
{b[46][0], b[46][1],b[46][2],b[46][3],b[46][4],b[46][5],b[46][6],b[46][7],b[46][8],b[46][9],b[46][10],b[46][11],b[46][12],b[46][13],b[46][14],b[46][15]} <= {b[45][0], b[45][1],b[45][2],b[45][3],b[45][4],b[45][5],b[45][6],b[45][7],b[45][8],b[45][9],b[45][10],b[45][11],b[45][12],b[45][13],b[45][14],b[45][15]}; 
{b[47][0], b[47][1],b[47][2],b[47][3],b[47][4],b[47][5],b[47][6],b[47][7],b[47][8],b[47][9],b[47][10],b[47][11],b[47][12],b[47][13],b[47][14],b[47][15]} <= {b[46][0], b[46][1],b[46][2],b[46][3],b[46][4],b[46][5],b[46][6],b[46][7],b[46][8],b[46][9],b[46][10],b[46][11],b[46][12],b[46][13],b[46][14],b[46][15]}; 
{b[48][0], b[48][1],b[48][2],b[48][3],b[48][4],b[48][5],b[48][6],b[48][7],b[48][8],b[48][9],b[48][10],b[48][11],b[48][12],b[48][13],b[48][14],b[48][15]} <= {b[47][0], b[47][1],b[47][2],b[47][3],b[47][4],b[47][5],b[47][6],b[47][7],b[47][8],b[47][9],b[47][10],b[47][11],b[47][12],b[47][13],b[47][14],b[47][15]}; 
{b[49][0], b[49][1],b[49][2],b[49][3],b[49][4],b[49][5],b[49][6],b[49][7],b[49][8],b[49][9],b[49][10],b[49][11],b[49][12],b[49][13],b[49][14],b[49][15]} <= {b[48][0], b[48][1],b[48][2],b[48][3],b[48][4],b[48][5],b[48][6],b[48][7],b[48][8],b[48][9],b[48][10],b[48][11],b[48][12],b[48][13],b[48][14],b[48][15]}; 
{b[50][0], b[50][1],b[50][2],b[50][3],b[50][4],b[50][5],b[50][6],b[50][7],b[50][8],b[50][9],b[50][10],b[50][11],b[50][12],b[50][13],b[50][14],b[50][15]} <= {b[49][0], b[49][1],b[49][2],b[49][3],b[49][4],b[49][5],b[49][6],b[49][7],b[49][8],b[49][9],b[49][10],b[49][11],b[49][12],b[49][13],b[49][14],b[49][15]}; 
{b[51][0], b[51][1],b[51][2],b[51][3],b[51][4],b[51][5],b[51][6],b[51][7],b[51][8],b[51][9],b[51][10],b[51][11],b[51][12],b[51][13],b[51][14],b[51][15]} <= {b[50][0], b[50][1],b[50][2],b[50][3],b[50][4],b[50][5],b[50][6],b[50][7],b[50][8],b[50][9],b[50][10],b[50][11],b[50][12],b[50][13],b[50][14],b[50][15]}; 
{b[52][0], b[52][1],b[52][2],b[52][3],b[52][4],b[52][5],b[52][6],b[52][7],b[52][8],b[52][9],b[52][10],b[52][11],b[52][12],b[52][13],b[52][14],b[52][15]} <= {b[51][0], b[51][1],b[51][2],b[51][3],b[51][4],b[51][5],b[51][6],b[51][7],b[51][8],b[51][9],b[51][10],b[51][11],b[51][12],b[51][13],b[51][14],b[51][15]}; 
{b[53][0], b[53][1],b[53][2],b[53][3],b[53][4],b[53][5],b[53][6],b[53][7],b[53][8],b[53][9],b[53][10],b[53][11],b[53][12],b[53][13],b[53][14],b[53][15]} <= {b[52][0], b[52][1],b[52][2],b[52][3],b[52][4],b[52][5],b[52][6],b[52][7],b[52][8],b[52][9],b[52][10],b[52][11],b[52][12],b[52][13],b[52][14],b[52][15]}; 
{b[54][0], b[54][1],b[54][2],b[54][3],b[54][4],b[54][5],b[54][6],b[54][7],b[54][8],b[54][9],b[54][10],b[54][11],b[54][12],b[54][13],b[54][14],b[54][15]} <= {b[53][0], b[53][1],b[53][2],b[53][3],b[53][4],b[53][5],b[53][6],b[53][7],b[53][8],b[53][9],b[53][10],b[53][11],b[53][12],b[53][13],b[53][14],b[53][15]}; 
{b[55][0], b[55][1],b[55][2],b[55][3],b[55][4],b[55][5],b[55][6],b[55][7],b[55][8],b[55][9],b[55][10],b[55][11],b[55][12],b[55][13],b[55][14],b[55][15]} <= {b[54][0], b[54][1],b[54][2],b[54][3],b[54][4],b[54][5],b[54][6],b[54][7],b[54][8],b[54][9],b[54][10],b[54][11],b[54][12],b[54][13],b[54][14],b[54][15]}; 
{b[56][0], b[56][1],b[56][2],b[56][3],b[56][4],b[56][5],b[56][6],b[56][7],b[56][8],b[56][9],b[56][10],b[56][11],b[56][12],b[56][13],b[56][14],b[56][15]} <= {b[55][0], b[55][1],b[55][2],b[55][3],b[55][4],b[55][5],b[55][6],b[55][7],b[55][8],b[55][9],b[55][10],b[55][11],b[55][12],b[55][13],b[55][14],b[55][15]}; 
{b[57][0], b[57][1],b[57][2],b[57][3],b[57][4],b[57][5],b[57][6],b[57][7],b[57][8],b[57][9],b[57][10],b[57][11],b[57][12],b[57][13],b[57][14],b[57][15]} <= {b[56][0], b[56][1],b[56][2],b[56][3],b[56][4],b[56][5],b[56][6],b[56][7],b[56][8],b[56][9],b[56][10],b[56][11],b[56][12],b[56][13],b[56][14],b[56][15]}; 
{b[58][0], b[58][1],b[58][2],b[58][3],b[58][4],b[58][5],b[58][6],b[58][7],b[58][8],b[58][9],b[58][10],b[58][11],b[58][12],b[58][13],b[58][14],b[58][15]} <= {b[57][0], b[57][1],b[57][2],b[57][3],b[57][4],b[57][5],b[57][6],b[57][7],b[57][8],b[57][9],b[57][10],b[57][11],b[57][12],b[57][13],b[57][14],b[57][15]}; 
{b[59][0], b[59][1],b[59][2],b[59][3],b[59][4],b[59][5],b[59][6],b[59][7],b[59][8],b[59][9],b[59][10],b[59][11],b[59][12],b[59][13],b[59][14],b[59][15]} <= {b[58][0], b[58][1],b[58][2],b[58][3],b[58][4],b[58][5],b[58][6],b[58][7],b[58][8],b[58][9],b[58][10],b[58][11],b[58][12],b[58][13],b[58][14],b[58][15]}; 
{b[60][0], b[60][1],b[60][2],b[60][3],b[60][4],b[60][5],b[60][6],b[60][7],b[60][8],b[60][9],b[60][10],b[60][11],b[60][12],b[60][13],b[60][14],b[60][15]} <= {b[59][0], b[59][1],b[59][2],b[59][3],b[59][4],b[59][5],b[59][6],b[59][7],b[59][8],b[59][9],b[59][10],b[59][11],b[59][12],b[59][13],b[59][14],b[59][15]}; 
{b[61][0], b[61][1],b[61][2],b[61][3],b[61][4],b[61][5],b[61][6],b[61][7],b[61][8],b[61][9],b[61][10],b[61][11],b[61][12],b[61][13],b[61][14],b[61][15]} <= {b[60][0], b[60][1],b[60][2],b[60][3],b[60][4],b[60][5],b[60][6],b[60][7],b[60][8],b[60][9],b[60][10],b[60][11],b[60][12],b[60][13],b[60][14],b[60][15]}; 
{b[62][0], b[62][1],b[62][2],b[62][3],b[62][4],b[62][5],b[62][6],b[62][7],b[62][8],b[62][9],b[62][10],b[62][11],b[62][12],b[62][13],b[62][14],b[62][15]} <= {b[61][0], b[61][1],b[61][2],b[61][3],b[61][4],b[61][5],b[61][6],b[61][7],b[61][8],b[61][9],b[61][10],b[61][11],b[61][12],b[61][13],b[61][14],b[61][15]}; 
{b[63][0], b[63][1],b[63][2],b[63][3],b[63][4],b[63][5],b[63][6],b[63][7],b[63][8],b[63][9],b[63][10],b[63][11],b[63][12],b[63][13],b[63][14],b[63][15]} <= {b[62][0], b[62][1],b[62][2],b[62][3],b[62][4],b[62][5],b[62][6],b[62][7],b[62][8],b[62][9],b[62][10],b[62][11],b[62][12],b[62][13],b[62][14],b[62][15]}; 
{b[64][0], b[64][1],b[64][2],b[64][3],b[64][4],b[64][5],b[64][6],b[64][7],b[64][8],b[64][9],b[64][10],b[64][11],b[64][12],b[64][13],b[64][14],b[64][15]} <= {b[63][0], b[63][1],b[63][2],b[63][3],b[63][4],b[63][5],b[63][6],b[63][7],b[63][8],b[63][9],b[63][10],b[63][11],b[63][12],b[63][13],b[63][14],b[63][15]}; 
{b[65][0], b[65][1],b[65][2],b[65][3],b[65][4],b[65][5],b[65][6],b[65][7],b[65][8],b[65][9],b[65][10],b[65][11],b[65][12],b[65][13],b[65][14],b[65][15]} <= {b[64][0], b[64][1],b[64][2],b[64][3],b[64][4],b[64][5],b[64][6],b[64][7],b[64][8],b[64][9],b[64][10],b[64][11],b[64][12],b[64][13],b[64][14],b[64][15]}; 
{b[66][0], b[66][1],b[66][2],b[66][3],b[66][4],b[66][5],b[66][6],b[66][7],b[66][8],b[66][9],b[66][10],b[66][11],b[66][12],b[66][13],b[66][14],b[66][15]} <= {b[65][0], b[65][1],b[65][2],b[65][3],b[65][4],b[65][5],b[65][6],b[65][7],b[65][8],b[65][9],b[65][10],b[65][11],b[65][12],b[65][13],b[65][14],b[65][15]}; 
{b[67][0], b[67][1],b[67][2],b[67][3],b[67][4],b[67][5],b[67][6],b[67][7],b[67][8],b[67][9],b[67][10],b[67][11],b[67][12],b[67][13],b[67][14],b[67][15]} <= {b[66][0], b[66][1],b[66][2],b[66][3],b[66][4],b[66][5],b[66][6],b[66][7],b[66][8],b[66][9],b[66][10],b[66][11],b[66][12],b[66][13],b[66][14],b[66][15]}; 
{b[68][0], b[68][1],b[68][2],b[68][3],b[68][4],b[68][5],b[68][6],b[68][7],b[68][8],b[68][9],b[68][10],b[68][11],b[68][12],b[68][13],b[68][14],b[68][15]} <= {b[67][0], b[67][1],b[67][2],b[67][3],b[67][4],b[67][5],b[67][6],b[67][7],b[67][8],b[67][9],b[67][10],b[67][11],b[67][12],b[67][13],b[67][14],b[67][15]}; 
{b[69][0], b[69][1],b[69][2],b[69][3],b[69][4],b[69][5],b[69][6],b[69][7],b[69][8],b[69][9],b[69][10],b[69][11],b[69][12],b[69][13],b[69][14],b[69][15]} <= {b[68][0], b[68][1],b[68][2],b[68][3],b[68][4],b[68][5],b[68][6],b[68][7],b[68][8],b[68][9],b[68][10],b[68][11],b[68][12],b[68][13],b[68][14],b[68][15]}; 
{b[70][0], b[70][1],b[70][2],b[70][3],b[70][4],b[70][5],b[70][6],b[70][7],b[70][8],b[70][9],b[70][10],b[70][11],b[70][12],b[70][13],b[70][14],b[70][15]} <= {b[69][0], b[69][1],b[69][2],b[69][3],b[69][4],b[69][5],b[69][6],b[69][7],b[69][8],b[69][9],b[69][10],b[69][11],b[69][12],b[69][13],b[69][14],b[69][15]}; 
{b[71][0], b[71][1],b[71][2],b[71][3],b[71][4],b[71][5],b[71][6],b[71][7],b[71][8],b[71][9],b[71][10],b[71][11],b[71][12],b[71][13],b[71][14],b[71][15]} <= {b[70][0], b[70][1],b[70][2],b[70][3],b[70][4],b[70][5],b[70][6],b[70][7],b[70][8],b[70][9],b[70][10],b[70][11],b[70][12],b[70][13],b[70][14],b[70][15]}; 
{b[72][0], b[72][1],b[72][2],b[72][3],b[72][4],b[72][5],b[72][6],b[72][7],b[72][8],b[72][9],b[72][10],b[72][11],b[72][12],b[72][13],b[72][14],b[72][15]} <= {b[71][0], b[71][1],b[71][2],b[71][3],b[71][4],b[71][5],b[71][6],b[71][7],b[71][8],b[71][9],b[71][10],b[71][11],b[71][12],b[71][13],b[71][14],b[71][15]}; 
{b[73][0], b[73][1],b[73][2],b[73][3],b[73][4],b[73][5],b[73][6],b[73][7],b[73][8],b[73][9],b[73][10],b[73][11],b[73][12],b[73][13],b[73][14],b[73][15]} <= {b[72][0], b[72][1],b[72][2],b[72][3],b[72][4],b[72][5],b[72][6],b[72][7],b[72][8],b[72][9],b[72][10],b[72][11],b[72][12],b[72][13],b[72][14],b[72][15]}; 
{b[74][0], b[74][1],b[74][2],b[74][3],b[74][4],b[74][5],b[74][6],b[74][7],b[74][8],b[74][9],b[74][10],b[74][11],b[74][12],b[74][13],b[74][14],b[74][15]} <= {b[73][0], b[73][1],b[73][2],b[73][3],b[73][4],b[73][5],b[73][6],b[73][7],b[73][8],b[73][9],b[73][10],b[73][11],b[73][12],b[73][13],b[73][14],b[73][15]}; 
{b[75][0], b[75][1],b[75][2],b[75][3],b[75][4],b[75][5],b[75][6],b[75][7],b[75][8],b[75][9],b[75][10],b[75][11],b[75][12],b[75][13],b[75][14],b[75][15]} <= {b[74][0], b[74][1],b[74][2],b[74][3],b[74][4],b[74][5],b[74][6],b[74][7],b[74][8],b[74][9],b[74][10],b[74][11],b[74][12],b[74][13],b[74][14],b[74][15]}; 
{b[76][0], b[76][1],b[76][2],b[76][3],b[76][4],b[76][5],b[76][6],b[76][7],b[76][8],b[76][9],b[76][10],b[76][11],b[76][12],b[76][13],b[76][14],b[76][15]} <= {b[75][0], b[75][1],b[75][2],b[75][3],b[75][4],b[75][5],b[75][6],b[75][7],b[75][8],b[75][9],b[75][10],b[75][11],b[75][12],b[75][13],b[75][14],b[75][15]}; 
{b[77][0], b[77][1],b[77][2],b[77][3],b[77][4],b[77][5],b[77][6],b[77][7],b[77][8],b[77][9],b[77][10],b[77][11],b[77][12],b[77][13],b[77][14],b[77][15]} <= {b[76][0], b[76][1],b[76][2],b[76][3],b[76][4],b[76][5],b[76][6],b[76][7],b[76][8],b[76][9],b[76][10],b[76][11],b[76][12],b[76][13],b[76][14],b[76][15]}; 
{b[78][0], b[78][1],b[78][2],b[78][3],b[78][4],b[78][5],b[78][6],b[78][7],b[78][8],b[78][9],b[78][10],b[78][11],b[78][12],b[78][13],b[78][14],b[78][15]} <= {b[77][0], b[77][1],b[77][2],b[77][3],b[77][4],b[77][5],b[77][6],b[77][7],b[77][8],b[77][9],b[77][10],b[77][11],b[77][12],b[77][13],b[77][14],b[77][15]}; 
{b[79][0], b[79][1],b[79][2],b[79][3],b[79][4],b[79][5],b[79][6],b[79][7],b[79][8],b[79][9],b[79][10],b[79][11],b[79][12],b[79][13],b[79][14],b[79][15]} <= {b[78][0], b[78][1],b[78][2],b[78][3],b[78][4],b[78][5],b[78][6],b[78][7],b[78][8],b[78][9],b[78][10],b[78][11],b[78][12],b[78][13],b[78][14],b[78][15]}; 
{b[80][0], b[80][1],b[80][2],b[80][3],b[80][4],b[80][5],b[80][6],b[80][7],b[80][8],b[80][9],b[80][10],b[80][11],b[80][12],b[80][13],b[80][14],b[80][15]} <= {b[79][0], b[79][1],b[79][2],b[79][3],b[79][4],b[79][5],b[79][6],b[79][7],b[79][8],b[79][9],b[79][10],b[79][11],b[79][12],b[79][13],b[79][14],b[79][15]}; 
{b[81][0], b[81][1],b[81][2],b[81][3],b[81][4],b[81][5],b[81][6],b[81][7],b[81][8],b[81][9],b[81][10],b[81][11],b[81][12],b[81][13],b[81][14],b[81][15]} <= {b[80][0], b[80][1],b[80][2],b[80][3],b[80][4],b[80][5],b[80][6],b[80][7],b[80][8],b[80][9],b[80][10],b[80][11],b[80][12],b[80][13],b[80][14],b[80][15]}; 
{b[82][0], b[82][1],b[82][2],b[82][3],b[82][4],b[82][5],b[82][6],b[82][7],b[82][8],b[82][9],b[82][10],b[82][11],b[82][12],b[82][13],b[82][14],b[82][15]} <= {b[81][0], b[81][1],b[81][2],b[81][3],b[81][4],b[81][5],b[81][6],b[81][7],b[81][8],b[81][9],b[81][10],b[81][11],b[81][12],b[81][13],b[81][14],b[81][15]}; 
{b[83][0], b[83][1],b[83][2],b[83][3],b[83][4],b[83][5],b[83][6],b[83][7],b[83][8],b[83][9],b[83][10],b[83][11],b[83][12],b[83][13],b[83][14],b[83][15]} <= {b[82][0], b[82][1],b[82][2],b[82][3],b[82][4],b[82][5],b[82][6],b[82][7],b[82][8],b[82][9],b[82][10],b[82][11],b[82][12],b[82][13],b[82][14],b[82][15]}; 
{b[84][0], b[84][1],b[84][2],b[84][3],b[84][4],b[84][5],b[84][6],b[84][7],b[84][8],b[84][9],b[84][10],b[84][11],b[84][12],b[84][13],b[84][14],b[84][15]} <= {b[83][0], b[83][1],b[83][2],b[83][3],b[83][4],b[83][5],b[83][6],b[83][7],b[83][8],b[83][9],b[83][10],b[83][11],b[83][12],b[83][13],b[83][14],b[83][15]}; 
{b[85][0], b[85][1],b[85][2],b[85][3],b[85][4],b[85][5],b[85][6],b[85][7],b[85][8],b[85][9],b[85][10],b[85][11],b[85][12],b[85][13],b[85][14],b[85][15]} <= {b[84][0], b[84][1],b[84][2],b[84][3],b[84][4],b[84][5],b[84][6],b[84][7],b[84][8],b[84][9],b[84][10],b[84][11],b[84][12],b[84][13],b[84][14],b[84][15]}; 
{b[86][0], b[86][1],b[86][2],b[86][3],b[86][4],b[86][5],b[86][6],b[86][7],b[86][8],b[86][9],b[86][10],b[86][11],b[86][12],b[86][13],b[86][14],b[86][15]} <= {b[85][0], b[85][1],b[85][2],b[85][3],b[85][4],b[85][5],b[85][6],b[85][7],b[85][8],b[85][9],b[85][10],b[85][11],b[85][12],b[85][13],b[85][14],b[85][15]}; 
{b[87][0], b[87][1],b[87][2],b[87][3],b[87][4],b[87][5],b[87][6],b[87][7],b[87][8],b[87][9],b[87][10],b[87][11],b[87][12],b[87][13],b[87][14],b[87][15]} <= {b[86][0], b[86][1],b[86][2],b[86][3],b[86][4],b[86][5],b[86][6],b[86][7],b[86][8],b[86][9],b[86][10],b[86][11],b[86][12],b[86][13],b[86][14],b[86][15]}; 
{b[88][0], b[88][1],b[88][2],b[88][3],b[88][4],b[88][5],b[88][6],b[88][7],b[88][8],b[88][9],b[88][10],b[88][11],b[88][12],b[88][13],b[88][14],b[88][15]} <= {b[87][0], b[87][1],b[87][2],b[87][3],b[87][4],b[87][5],b[87][6],b[87][7],b[87][8],b[87][9],b[87][10],b[87][11],b[87][12],b[87][13],b[87][14],b[87][15]}; 
{b[89][0], b[89][1],b[89][2],b[89][3],b[89][4],b[89][5],b[89][6],b[89][7],b[89][8],b[89][9],b[89][10],b[89][11],b[89][12],b[89][13],b[89][14],b[89][15]} <= {b[88][0], b[88][1],b[88][2],b[88][3],b[88][4],b[88][5],b[88][6],b[88][7],b[88][8],b[88][9],b[88][10],b[88][11],b[88][12],b[88][13],b[88][14],b[88][15]}; 
{b[90][0], b[90][1],b[90][2],b[90][3],b[90][4],b[90][5],b[90][6],b[90][7],b[90][8],b[90][9],b[90][10],b[90][11],b[90][12],b[90][13],b[90][14],b[90][15]} <= {b[89][0], b[89][1],b[89][2],b[89][3],b[89][4],b[89][5],b[89][6],b[89][7],b[89][8],b[89][9],b[89][10],b[89][11],b[89][12],b[89][13],b[89][14],b[89][15]}; 
{b[91][0], b[91][1],b[91][2],b[91][3],b[91][4],b[91][5],b[91][6],b[91][7],b[91][8],b[91][9],b[91][10],b[91][11],b[91][12],b[91][13],b[91][14],b[91][15]} <= {b[90][0], b[90][1],b[90][2],b[90][3],b[90][4],b[90][5],b[90][6],b[90][7],b[90][8],b[90][9],b[90][10],b[90][11],b[90][12],b[90][13],b[90][14],b[90][15]}; 
{b[92][0], b[92][1],b[92][2],b[92][3],b[92][4],b[92][5],b[92][6],b[92][7],b[92][8],b[92][9],b[92][10],b[92][11],b[92][12],b[92][13],b[92][14],b[92][15]} <= {b[91][0], b[91][1],b[91][2],b[91][3],b[91][4],b[91][5],b[91][6],b[91][7],b[91][8],b[91][9],b[91][10],b[91][11],b[91][12],b[91][13],b[91][14],b[91][15]}; 
{b[93][0], b[93][1],b[93][2],b[93][3],b[93][4],b[93][5],b[93][6],b[93][7],b[93][8],b[93][9],b[93][10],b[93][11],b[93][12],b[93][13],b[93][14],b[93][15]} <= {b[92][0], b[92][1],b[92][2],b[92][3],b[92][4],b[92][5],b[92][6],b[92][7],b[92][8],b[92][9],b[92][10],b[92][11],b[92][12],b[92][13],b[92][14],b[92][15]}; 
{b[94][0], b[94][1],b[94][2],b[94][3],b[94][4],b[94][5],b[94][6],b[94][7],b[94][8],b[94][9],b[94][10],b[94][11],b[94][12],b[94][13],b[94][14],b[94][15]} <= {b[93][0], b[93][1],b[93][2],b[93][3],b[93][4],b[93][5],b[93][6],b[93][7],b[93][8],b[93][9],b[93][10],b[93][11],b[93][12],b[93][13],b[93][14],b[93][15]}; 
{b[95][0], b[95][1],b[95][2],b[95][3],b[95][4],b[95][5],b[95][6],b[95][7],b[95][8],b[95][9],b[95][10],b[95][11],b[95][12],b[95][13],b[95][14],b[95][15]} <= {b[94][0], b[94][1],b[94][2],b[94][3],b[94][4],b[94][5],b[94][6],b[94][7],b[94][8],b[94][9],b[94][10],b[94][11],b[94][12],b[94][13],b[94][14],b[94][15]}; 
{b[96][0], b[96][1],b[96][2],b[96][3],b[96][4],b[96][5],b[96][6],b[96][7],b[96][8],b[96][9],b[96][10],b[96][11],b[96][12],b[96][13],b[96][14],b[96][15]} <= {b[95][0], b[95][1],b[95][2],b[95][3],b[95][4],b[95][5],b[95][6],b[95][7],b[95][8],b[95][9],b[95][10],b[95][11],b[95][12],b[95][13],b[95][14],b[95][15]}; 
{b[97][0], b[97][1],b[97][2],b[97][3],b[97][4],b[97][5],b[97][6],b[97][7],b[97][8],b[97][9],b[97][10],b[97][11],b[97][12],b[97][13],b[97][14],b[97][15]} <= {b[96][0], b[96][1],b[96][2],b[96][3],b[96][4],b[96][5],b[96][6],b[96][7],b[96][8],b[96][9],b[96][10],b[96][11],b[96][12],b[96][13],b[96][14],b[96][15]}; 
{b[98][0], b[98][1],b[98][2],b[98][3],b[98][4],b[98][5],b[98][6],b[98][7],b[98][8],b[98][9],b[98][10],b[98][11],b[98][12],b[98][13],b[98][14],b[98][15]} <= {b[97][0], b[97][1],b[97][2],b[97][3],b[97][4],b[97][5],b[97][6],b[97][7],b[97][8],b[97][9],b[97][10],b[97][11],b[97][12],b[97][13],b[97][14],b[97][15]}; 
{b[99][0], b[99][1],b[99][2],b[99][3],b[99][4],b[99][5],b[99][6],b[99][7],b[99][8],b[99][9],b[99][10],b[99][11],b[99][12],b[99][13],b[99][14],b[99][15]} <= {b[98][0], b[98][1],b[98][2],b[98][3],b[98][4],b[98][5],b[98][6],b[98][7],b[98][8],b[98][9],b[98][10],b[98][11],b[98][12],b[98][13],b[98][14],b[98][15]}; 
{b[100][0], b[100][1],b[100][2],b[100][3],b[100][4],b[100][5],b[100][6],b[100][7],b[100][8],b[100][9],b[100][10],b[100][11],b[100][12],b[100][13],b[100][14],b[100][15]} <= {b[99][0], b[99][1],b[99][2],b[99][3],b[99][4],b[99][5],b[99][6],b[99][7],b[99][8],b[99][9],b[99][10],b[99][11],b[99][12],b[99][13],b[99][14],b[99][15]}; 
{b[101][0], b[101][1],b[101][2],b[101][3],b[101][4],b[101][5],b[101][6],b[101][7],b[101][8],b[101][9],b[101][10],b[101][11],b[101][12],b[101][13],b[101][14],b[101][15]} <= {b[100][0], b[100][1],b[100][2],b[100][3],b[100][4],b[100][5],b[100][6],b[100][7],b[100][8],b[100][9],b[100][10],b[100][11],b[100][12],b[100][13],b[100][14],b[100][15]}; 
{b[102][0], b[102][1],b[102][2],b[102][3],b[102][4],b[102][5],b[102][6],b[102][7],b[102][8],b[102][9],b[102][10],b[102][11],b[102][12],b[102][13],b[102][14],b[102][15]} <= {b[101][0], b[101][1],b[101][2],b[101][3],b[101][4],b[101][5],b[101][6],b[101][7],b[101][8],b[101][9],b[101][10],b[101][11],b[101][12],b[101][13],b[101][14],b[101][15]}; 
{b[103][0], b[103][1],b[103][2],b[103][3],b[103][4],b[103][5],b[103][6],b[103][7],b[103][8],b[103][9],b[103][10],b[103][11],b[103][12],b[103][13],b[103][14],b[103][15]} <= {b[102][0], b[102][1],b[102][2],b[102][3],b[102][4],b[102][5],b[102][6],b[102][7],b[102][8],b[102][9],b[102][10],b[102][11],b[102][12],b[102][13],b[102][14],b[102][15]}; 
{b[104][0], b[104][1],b[104][2],b[104][3],b[104][4],b[104][5],b[104][6],b[104][7],b[104][8],b[104][9],b[104][10],b[104][11],b[104][12],b[104][13],b[104][14],b[104][15]} <= {b[103][0], b[103][1],b[103][2],b[103][3],b[103][4],b[103][5],b[103][6],b[103][7],b[103][8],b[103][9],b[103][10],b[103][11],b[103][12],b[103][13],b[103][14],b[103][15]}; 
{b[105][0], b[105][1],b[105][2],b[105][3],b[105][4],b[105][5],b[105][6],b[105][7],b[105][8],b[105][9],b[105][10],b[105][11],b[105][12],b[105][13],b[105][14],b[105][15]} <= {b[104][0], b[104][1],b[104][2],b[104][3],b[104][4],b[104][5],b[104][6],b[104][7],b[104][8],b[104][9],b[104][10],b[104][11],b[104][12],b[104][13],b[104][14],b[104][15]}; 
{b[106][0], b[106][1],b[106][2],b[106][3],b[106][4],b[106][5],b[106][6],b[106][7],b[106][8],b[106][9],b[106][10],b[106][11],b[106][12],b[106][13],b[106][14],b[106][15]} <= {b[105][0], b[105][1],b[105][2],b[105][3],b[105][4],b[105][5],b[105][6],b[105][7],b[105][8],b[105][9],b[105][10],b[105][11],b[105][12],b[105][13],b[105][14],b[105][15]}; 
{b[107][0], b[107][1],b[107][2],b[107][3],b[107][4],b[107][5],b[107][6],b[107][7],b[107][8],b[107][9],b[107][10],b[107][11],b[107][12],b[107][13],b[107][14],b[107][15]} <= {b[106][0], b[106][1],b[106][2],b[106][3],b[106][4],b[106][5],b[106][6],b[106][7],b[106][8],b[106][9],b[106][10],b[106][11],b[106][12],b[106][13],b[106][14],b[106][15]}; 
{b[108][0], b[108][1],b[108][2],b[108][3],b[108][4],b[108][5],b[108][6],b[108][7],b[108][8],b[108][9],b[108][10],b[108][11],b[108][12],b[108][13],b[108][14],b[108][15]} <= {b[107][0], b[107][1],b[107][2],b[107][3],b[107][4],b[107][5],b[107][6],b[107][7],b[107][8],b[107][9],b[107][10],b[107][11],b[107][12],b[107][13],b[107][14],b[107][15]}; 
{b[109][0], b[109][1],b[109][2],b[109][3],b[109][4],b[109][5],b[109][6],b[109][7],b[109][8],b[109][9],b[109][10],b[109][11],b[109][12],b[109][13],b[109][14],b[109][15]} <= {b[108][0], b[108][1],b[108][2],b[108][3],b[108][4],b[108][5],b[108][6],b[108][7],b[108][8],b[108][9],b[108][10],b[108][11],b[108][12],b[108][13],b[108][14],b[108][15]}; 
{b[110][0], b[110][1],b[110][2],b[110][3],b[110][4],b[110][5],b[110][6],b[110][7],b[110][8],b[110][9],b[110][10],b[110][11],b[110][12],b[110][13],b[110][14],b[110][15]} <= {b[109][0], b[109][1],b[109][2],b[109][3],b[109][4],b[109][5],b[109][6],b[109][7],b[109][8],b[109][9],b[109][10],b[109][11],b[109][12],b[109][13],b[109][14],b[109][15]}; 
{b[111][0], b[111][1],b[111][2],b[111][3],b[111][4],b[111][5],b[111][6],b[111][7],b[111][8],b[111][9],b[111][10],b[111][11],b[111][12],b[111][13],b[111][14],b[111][15]} <= {b[110][0], b[110][1],b[110][2],b[110][3],b[110][4],b[110][5],b[110][6],b[110][7],b[110][8],b[110][9],b[110][10],b[110][11],b[110][12],b[110][13],b[110][14],b[110][15]}; 
{b[112][0], b[112][1],b[112][2],b[112][3],b[112][4],b[112][5],b[112][6],b[112][7],b[112][8],b[112][9],b[112][10],b[112][11],b[112][12],b[112][13],b[112][14],b[112][15]} <= {b[111][0], b[111][1],b[111][2],b[111][3],b[111][4],b[111][5],b[111][6],b[111][7],b[111][8],b[111][9],b[111][10],b[111][11],b[111][12],b[111][13],b[111][14],b[111][15]}; 
{b[113][0], b[113][1],b[113][2],b[113][3],b[113][4],b[113][5],b[113][6],b[113][7],b[113][8],b[113][9],b[113][10],b[113][11],b[113][12],b[113][13],b[113][14],b[113][15]} <= {b[112][0], b[112][1],b[112][2],b[112][3],b[112][4],b[112][5],b[112][6],b[112][7],b[112][8],b[112][9],b[112][10],b[112][11],b[112][12],b[112][13],b[112][14],b[112][15]}; 
{b[114][0], b[114][1],b[114][2],b[114][3],b[114][4],b[114][5],b[114][6],b[114][7],b[114][8],b[114][9],b[114][10],b[114][11],b[114][12],b[114][13],b[114][14],b[114][15]} <= {b[113][0], b[113][1],b[113][2],b[113][3],b[113][4],b[113][5],b[113][6],b[113][7],b[113][8],b[113][9],b[113][10],b[113][11],b[113][12],b[113][13],b[113][14],b[113][15]}; 
{b[115][0], b[115][1],b[115][2],b[115][3],b[115][4],b[115][5],b[115][6],b[115][7],b[115][8],b[115][9],b[115][10],b[115][11],b[115][12],b[115][13],b[115][14],b[115][15]} <= {b[114][0], b[114][1],b[114][2],b[114][3],b[114][4],b[114][5],b[114][6],b[114][7],b[114][8],b[114][9],b[114][10],b[114][11],b[114][12],b[114][13],b[114][14],b[114][15]}; 
{b[116][0], b[116][1],b[116][2],b[116][3],b[116][4],b[116][5],b[116][6],b[116][7],b[116][8],b[116][9],b[116][10],b[116][11],b[116][12],b[116][13],b[116][14],b[116][15]} <= {b[115][0], b[115][1],b[115][2],b[115][3],b[115][4],b[115][5],b[115][6],b[115][7],b[115][8],b[115][9],b[115][10],b[115][11],b[115][12],b[115][13],b[115][14],b[115][15]}; 
{b[117][0], b[117][1],b[117][2],b[117][3],b[117][4],b[117][5],b[117][6],b[117][7],b[117][8],b[117][9],b[117][10],b[117][11],b[117][12],b[117][13],b[117][14],b[117][15]} <= {b[116][0], b[116][1],b[116][2],b[116][3],b[116][4],b[116][5],b[116][6],b[116][7],b[116][8],b[116][9],b[116][10],b[116][11],b[116][12],b[116][13],b[116][14],b[116][15]}; 
{b[118][0], b[118][1],b[118][2],b[118][3],b[118][4],b[118][5],b[118][6],b[118][7],b[118][8],b[118][9],b[118][10],b[118][11],b[118][12],b[118][13],b[118][14],b[118][15]} <= {b[117][0], b[117][1],b[117][2],b[117][3],b[117][4],b[117][5],b[117][6],b[117][7],b[117][8],b[117][9],b[117][10],b[117][11],b[117][12],b[117][13],b[117][14],b[117][15]}; 
{b[119][0], b[119][1],b[119][2],b[119][3],b[119][4],b[119][5],b[119][6],b[119][7],b[119][8],b[119][9],b[119][10],b[119][11],b[119][12],b[119][13],b[119][14],b[119][15]} <= {b[118][0], b[118][1],b[118][2],b[118][3],b[118][4],b[118][5],b[118][6],b[118][7],b[118][8],b[118][9],b[118][10],b[118][11],b[118][12],b[118][13],b[118][14],b[118][15]}; 
{b[120][0], b[120][1],b[120][2],b[120][3],b[120][4],b[120][5],b[120][6],b[120][7],b[120][8],b[120][9],b[120][10],b[120][11],b[120][12],b[120][13],b[120][14],b[120][15]} <= {b[119][0], b[119][1],b[119][2],b[119][3],b[119][4],b[119][5],b[119][6],b[119][7],b[119][8],b[119][9],b[119][10],b[119][11],b[119][12],b[119][13],b[119][14],b[119][15]}; 
{b[121][0], b[121][1],b[121][2],b[121][3],b[121][4],b[121][5],b[121][6],b[121][7],b[121][8],b[121][9],b[121][10],b[121][11],b[121][12],b[121][13],b[121][14],b[121][15]} <= {b[120][0], b[120][1],b[120][2],b[120][3],b[120][4],b[120][5],b[120][6],b[120][7],b[120][8],b[120][9],b[120][10],b[120][11],b[120][12],b[120][13],b[120][14],b[120][15]}; 
{b[122][0], b[122][1],b[122][2],b[122][3],b[122][4],b[122][5],b[122][6],b[122][7],b[122][8],b[122][9],b[122][10],b[122][11],b[122][12],b[122][13],b[122][14],b[122][15]} <= {b[121][0], b[121][1],b[121][2],b[121][3],b[121][4],b[121][5],b[121][6],b[121][7],b[121][8],b[121][9],b[121][10],b[121][11],b[121][12],b[121][13],b[121][14],b[121][15]}; 
{b[123][0], b[123][1],b[123][2],b[123][3],b[123][4],b[123][5],b[123][6],b[123][7],b[123][8],b[123][9],b[123][10],b[123][11],b[123][12],b[123][13],b[123][14],b[123][15]} <= {b[122][0], b[122][1],b[122][2],b[122][3],b[122][4],b[122][5],b[122][6],b[122][7],b[122][8],b[122][9],b[122][10],b[122][11],b[122][12],b[122][13],b[122][14],b[122][15]}; 
{b[124][0], b[124][1],b[124][2],b[124][3],b[124][4],b[124][5],b[124][6],b[124][7],b[124][8],b[124][9],b[124][10],b[124][11],b[124][12],b[124][13],b[124][14],b[124][15]} <= {b[123][0], b[123][1],b[123][2],b[123][3],b[123][4],b[123][5],b[123][6],b[123][7],b[123][8],b[123][9],b[123][10],b[123][11],b[123][12],b[123][13],b[123][14],b[123][15]}; 
{b[125][0], b[125][1],b[125][2],b[125][3],b[125][4],b[125][5],b[125][6],b[125][7],b[125][8],b[125][9],b[125][10],b[125][11],b[125][12],b[125][13],b[125][14],b[125][15]} <= {b[124][0], b[124][1],b[124][2],b[124][3],b[124][4],b[124][5],b[124][6],b[124][7],b[124][8],b[124][9],b[124][10],b[124][11],b[124][12],b[124][13],b[124][14],b[124][15]}; 
{b[126][0], b[126][1],b[126][2],b[126][3],b[126][4],b[126][5],b[126][6],b[126][7],b[126][8],b[126][9],b[126][10],b[126][11],b[126][12],b[126][13],b[126][14],b[126][15]} <= {b[125][0], b[125][1],b[125][2],b[125][3],b[125][4],b[125][5],b[125][6],b[125][7],b[125][8],b[125][9],b[125][10],b[125][11],b[125][12],b[125][13],b[125][14],b[125][15]}; 
{b[127][0], b[127][1],b[127][2],b[127][3],b[127][4],b[127][5],b[127][6],b[127][7],b[127][8],b[127][9],b[127][10],b[127][11],b[127][12],b[127][13],b[127][14],b[127][15]} <= {b[126][0], b[126][1],b[126][2],b[126][3],b[126][4],b[126][5],b[126][6],b[126][7],b[126][8],b[126][9],b[126][10],b[126][11],b[126][12],b[126][13],b[126][14],b[126][15]}; 
{b[128][0], b[128][1],b[128][2],b[128][3],b[128][4],b[128][5],b[128][6],b[128][7],b[128][8],b[128][9],b[128][10],b[128][11],b[128][12],b[128][13],b[128][14],b[128][15]} <= {b[127][0], b[127][1],b[127][2],b[127][3],b[127][4],b[127][5],b[127][6],b[127][7],b[127][8],b[127][9],b[127][10],b[127][11],b[127][12],b[127][13],b[127][14],b[127][15]}; 
{b[129][0], b[129][1],b[129][2],b[129][3],b[129][4],b[129][5],b[129][6],b[129][7],b[129][8],b[129][9],b[129][10],b[129][11],b[129][12],b[129][13],b[129][14],b[129][15]} <= {b[128][0], b[128][1],b[128][2],b[128][3],b[128][4],b[128][5],b[128][6],b[128][7],b[128][8],b[128][9],b[128][10],b[128][11],b[128][12],b[128][13],b[128][14],b[128][15]}; 
{b[130][0], b[130][1],b[130][2],b[130][3],b[130][4],b[130][5],b[130][6],b[130][7],b[130][8],b[130][9],b[130][10],b[130][11],b[130][12],b[130][13],b[130][14],b[130][15]} <= {b[129][0], b[129][1],b[129][2],b[129][3],b[129][4],b[129][5],b[129][6],b[129][7],b[129][8],b[129][9],b[129][10],b[129][11],b[129][12],b[129][13],b[129][14],b[129][15]}; 
{b[131][0], b[131][1],b[131][2],b[131][3],b[131][4],b[131][5],b[131][6],b[131][7],b[131][8],b[131][9],b[131][10],b[131][11],b[131][12],b[131][13],b[131][14],b[131][15]} <= {b[130][0], b[130][1],b[130][2],b[130][3],b[130][4],b[130][5],b[130][6],b[130][7],b[130][8],b[130][9],b[130][10],b[130][11],b[130][12],b[130][13],b[130][14],b[130][15]}; 
{b[132][0], b[132][1],b[132][2],b[132][3],b[132][4],b[132][5],b[132][6],b[132][7],b[132][8],b[132][9],b[132][10],b[132][11],b[132][12],b[132][13],b[132][14],b[132][15]} <= {b[131][0], b[131][1],b[131][2],b[131][3],b[131][4],b[131][5],b[131][6],b[131][7],b[131][8],b[131][9],b[131][10],b[131][11],b[131][12],b[131][13],b[131][14],b[131][15]}; 
{b[133][0], b[133][1],b[133][2],b[133][3],b[133][4],b[133][5],b[133][6],b[133][7],b[133][8],b[133][9],b[133][10],b[133][11],b[133][12],b[133][13],b[133][14],b[133][15]} <= {b[132][0], b[132][1],b[132][2],b[132][3],b[132][4],b[132][5],b[132][6],b[132][7],b[132][8],b[132][9],b[132][10],b[132][11],b[132][12],b[132][13],b[132][14],b[132][15]}; 
{b[134][0], b[134][1],b[134][2],b[134][3],b[134][4],b[134][5],b[134][6],b[134][7],b[134][8],b[134][9],b[134][10],b[134][11],b[134][12],b[134][13],b[134][14],b[134][15]} <= {b[133][0], b[133][1],b[133][2],b[133][3],b[133][4],b[133][5],b[133][6],b[133][7],b[133][8],b[133][9],b[133][10],b[133][11],b[133][12],b[133][13],b[133][14],b[133][15]}; 
{b[135][0], b[135][1],b[135][2],b[135][3],b[135][4],b[135][5],b[135][6],b[135][7],b[135][8],b[135][9],b[135][10],b[135][11],b[135][12],b[135][13],b[135][14],b[135][15]} <= {b[134][0], b[134][1],b[134][2],b[134][3],b[134][4],b[134][5],b[134][6],b[134][7],b[134][8],b[134][9],b[134][10],b[134][11],b[134][12],b[134][13],b[134][14],b[134][15]}; 
{b[136][0], b[136][1],b[136][2],b[136][3],b[136][4],b[136][5],b[136][6],b[136][7],b[136][8],b[136][9],b[136][10],b[136][11],b[136][12],b[136][13],b[136][14],b[136][15]} <= {b[135][0], b[135][1],b[135][2],b[135][3],b[135][4],b[135][5],b[135][6],b[135][7],b[135][8],b[135][9],b[135][10],b[135][11],b[135][12],b[135][13],b[135][14],b[135][15]}; 
{b[137][0], b[137][1],b[137][2],b[137][3],b[137][4],b[137][5],b[137][6],b[137][7],b[137][8],b[137][9],b[137][10],b[137][11],b[137][12],b[137][13],b[137][14],b[137][15]} <= {b[136][0], b[136][1],b[136][2],b[136][3],b[136][4],b[136][5],b[136][6],b[136][7],b[136][8],b[136][9],b[136][10],b[136][11],b[136][12],b[136][13],b[136][14],b[136][15]}; 
{b[138][0], b[138][1],b[138][2],b[138][3],b[138][4],b[138][5],b[138][6],b[138][7],b[138][8],b[138][9],b[138][10],b[138][11],b[138][12],b[138][13],b[138][14],b[138][15]} <= {b[137][0], b[137][1],b[137][2],b[137][3],b[137][4],b[137][5],b[137][6],b[137][7],b[137][8],b[137][9],b[137][10],b[137][11],b[137][12],b[137][13],b[137][14],b[137][15]}; 
{b[139][0], b[139][1],b[139][2],b[139][3],b[139][4],b[139][5],b[139][6],b[139][7],b[139][8],b[139][9],b[139][10],b[139][11],b[139][12],b[139][13],b[139][14],b[139][15]} <= {b[138][0], b[138][1],b[138][2],b[138][3],b[138][4],b[138][5],b[138][6],b[138][7],b[138][8],b[138][9],b[138][10],b[138][11],b[138][12],b[138][13],b[138][14],b[138][15]}; 
{b[140][0], b[140][1],b[140][2],b[140][3],b[140][4],b[140][5],b[140][6],b[140][7],b[140][8],b[140][9],b[140][10],b[140][11],b[140][12],b[140][13],b[140][14],b[140][15]} <= {b[139][0], b[139][1],b[139][2],b[139][3],b[139][4],b[139][5],b[139][6],b[139][7],b[139][8],b[139][9],b[139][10],b[139][11],b[139][12],b[139][13],b[139][14],b[139][15]}; 
{b[141][0], b[141][1],b[141][2],b[141][3],b[141][4],b[141][5],b[141][6],b[141][7],b[141][8],b[141][9],b[141][10],b[141][11],b[141][12],b[141][13],b[141][14],b[141][15]} <= {b[140][0], b[140][1],b[140][2],b[140][3],b[140][4],b[140][5],b[140][6],b[140][7],b[140][8],b[140][9],b[140][10],b[140][11],b[140][12],b[140][13],b[140][14],b[140][15]}; 
{b[142][0], b[142][1],b[142][2],b[142][3],b[142][4],b[142][5],b[142][6],b[142][7],b[142][8],b[142][9],b[142][10],b[142][11],b[142][12],b[142][13],b[142][14],b[142][15]} <= {b[141][0], b[141][1],b[141][2],b[141][3],b[141][4],b[141][5],b[141][6],b[141][7],b[141][8],b[141][9],b[141][10],b[141][11],b[141][12],b[141][13],b[141][14],b[141][15]}; 
{b[143][0], b[143][1],b[143][2],b[143][3],b[143][4],b[143][5],b[143][6],b[143][7],b[143][8],b[143][9],b[143][10],b[143][11],b[143][12],b[143][13],b[143][14],b[143][15]} <= {b[142][0], b[142][1],b[142][2],b[142][3],b[142][4],b[142][5],b[142][6],b[142][7],b[142][8],b[142][9],b[142][10],b[142][11],b[142][12],b[142][13],b[142][14],b[142][15]}; 
{b[144][0], b[144][1],b[144][2],b[144][3],b[144][4],b[144][5],b[144][6],b[144][7],b[144][8],b[144][9],b[144][10],b[144][11],b[144][12],b[144][13],b[144][14],b[144][15]} <= {b[143][0], b[143][1],b[143][2],b[143][3],b[143][4],b[143][5],b[143][6],b[143][7],b[143][8],b[143][9],b[143][10],b[143][11],b[143][12],b[143][13],b[143][14],b[143][15]}; 
{b[145][0], b[145][1],b[145][2],b[145][3],b[145][4],b[145][5],b[145][6],b[145][7],b[145][8],b[145][9],b[145][10],b[145][11],b[145][12],b[145][13],b[145][14],b[145][15]} <= {b[144][0], b[144][1],b[144][2],b[144][3],b[144][4],b[144][5],b[144][6],b[144][7],b[144][8],b[144][9],b[144][10],b[144][11],b[144][12],b[144][13],b[144][14],b[144][15]}; 
{b[146][0], b[146][1],b[146][2],b[146][3],b[146][4],b[146][5],b[146][6],b[146][7],b[146][8],b[146][9],b[146][10],b[146][11],b[146][12],b[146][13],b[146][14],b[146][15]} <= {b[145][0], b[145][1],b[145][2],b[145][3],b[145][4],b[145][5],b[145][6],b[145][7],b[145][8],b[145][9],b[145][10],b[145][11],b[145][12],b[145][13],b[145][14],b[145][15]}; 
{b[147][0], b[147][1],b[147][2],b[147][3],b[147][4],b[147][5],b[147][6],b[147][7],b[147][8],b[147][9],b[147][10],b[147][11],b[147][12],b[147][13],b[147][14],b[147][15]} <= {b[146][0], b[146][1],b[146][2],b[146][3],b[146][4],b[146][5],b[146][6],b[146][7],b[146][8],b[146][9],b[146][10],b[146][11],b[146][12],b[146][13],b[146][14],b[146][15]}; 
{b[148][0], b[148][1],b[148][2],b[148][3],b[148][4],b[148][5],b[148][6],b[148][7],b[148][8],b[148][9],b[148][10],b[148][11],b[148][12],b[148][13],b[148][14],b[148][15]} <= {b[147][0], b[147][1],b[147][2],b[147][3],b[147][4],b[147][5],b[147][6],b[147][7],b[147][8],b[147][9],b[147][10],b[147][11],b[147][12],b[147][13],b[147][14],b[147][15]}; 
{b[149][0], b[149][1],b[149][2],b[149][3],b[149][4],b[149][5],b[149][6],b[149][7],b[149][8],b[149][9],b[149][10],b[149][11],b[149][12],b[149][13],b[149][14],b[149][15]} <= {b[148][0], b[148][1],b[148][2],b[148][3],b[148][4],b[148][5],b[148][6],b[148][7],b[148][8],b[148][9],b[148][10],b[148][11],b[148][12],b[148][13],b[148][14],b[148][15]}; 
{b[150][0], b[150][1],b[150][2],b[150][3],b[150][4],b[150][5],b[150][6],b[150][7],b[150][8],b[150][9],b[150][10],b[150][11],b[150][12],b[150][13],b[150][14],b[150][15]} <= {b[149][0], b[149][1],b[149][2],b[149][3],b[149][4],b[149][5],b[149][6],b[149][7],b[149][8],b[149][9],b[149][10],b[149][11],b[149][12],b[149][13],b[149][14],b[149][15]}; 
{b[151][0], b[151][1],b[151][2],b[151][3],b[151][4],b[151][5],b[151][6],b[151][7],b[151][8],b[151][9],b[151][10],b[151][11],b[151][12],b[151][13],b[151][14],b[151][15]} <= {b[150][0], b[150][1],b[150][2],b[150][3],b[150][4],b[150][5],b[150][6],b[150][7],b[150][8],b[150][9],b[150][10],b[150][11],b[150][12],b[150][13],b[150][14],b[150][15]}; 
{b[152][0], b[152][1],b[152][2],b[152][3],b[152][4],b[152][5],b[152][6],b[152][7],b[152][8],b[152][9],b[152][10],b[152][11],b[152][12],b[152][13],b[152][14],b[152][15]} <= {b[151][0], b[151][1],b[151][2],b[151][3],b[151][4],b[151][5],b[151][6],b[151][7],b[151][8],b[151][9],b[151][10],b[151][11],b[151][12],b[151][13],b[151][14],b[151][15]}; 
{b[153][0], b[153][1],b[153][2],b[153][3],b[153][4],b[153][5],b[153][6],b[153][7],b[153][8],b[153][9],b[153][10],b[153][11],b[153][12],b[153][13],b[153][14],b[153][15]} <= {b[152][0], b[152][1],b[152][2],b[152][3],b[152][4],b[152][5],b[152][6],b[152][7],b[152][8],b[152][9],b[152][10],b[152][11],b[152][12],b[152][13],b[152][14],b[152][15]}; 
{b[154][0], b[154][1],b[154][2],b[154][3],b[154][4],b[154][5],b[154][6],b[154][7],b[154][8],b[154][9],b[154][10],b[154][11],b[154][12],b[154][13],b[154][14],b[154][15]} <= {b[153][0], b[153][1],b[153][2],b[153][3],b[153][4],b[153][5],b[153][6],b[153][7],b[153][8],b[153][9],b[153][10],b[153][11],b[153][12],b[153][13],b[153][14],b[153][15]}; 
{b[155][0], b[155][1],b[155][2],b[155][3],b[155][4],b[155][5],b[155][6],b[155][7],b[155][8],b[155][9],b[155][10],b[155][11],b[155][12],b[155][13],b[155][14],b[155][15]} <= {b[154][0], b[154][1],b[154][2],b[154][3],b[154][4],b[154][5],b[154][6],b[154][7],b[154][8],b[154][9],b[154][10],b[154][11],b[154][12],b[154][13],b[154][14],b[154][15]}; 
{b[156][0], b[156][1],b[156][2],b[156][3],b[156][4],b[156][5],b[156][6],b[156][7],b[156][8],b[156][9],b[156][10],b[156][11],b[156][12],b[156][13],b[156][14],b[156][15]} <= {b[155][0], b[155][1],b[155][2],b[155][3],b[155][4],b[155][5],b[155][6],b[155][7],b[155][8],b[155][9],b[155][10],b[155][11],b[155][12],b[155][13],b[155][14],b[155][15]}; 
{b[157][0], b[157][1],b[157][2],b[157][3],b[157][4],b[157][5],b[157][6],b[157][7],b[157][8],b[157][9],b[157][10],b[157][11],b[157][12],b[157][13],b[157][14],b[157][15]} <= {b[156][0], b[156][1],b[156][2],b[156][3],b[156][4],b[156][5],b[156][6],b[156][7],b[156][8],b[156][9],b[156][10],b[156][11],b[156][12],b[156][13],b[156][14],b[156][15]}; 
{b[158][0], b[158][1],b[158][2],b[158][3],b[158][4],b[158][5],b[158][6],b[158][7],b[158][8],b[158][9],b[158][10],b[158][11],b[158][12],b[158][13],b[158][14],b[158][15]} <= {b[157][0], b[157][1],b[157][2],b[157][3],b[157][4],b[157][5],b[157][6],b[157][7],b[157][8],b[157][9],b[157][10],b[157][11],b[157][12],b[157][13],b[157][14],b[157][15]}; 
{b[159][0], b[159][1],b[159][2],b[159][3],b[159][4],b[159][5],b[159][6],b[159][7],b[159][8],b[159][9],b[159][10],b[159][11],b[159][12],b[159][13],b[159][14],b[159][15]} <= {b[158][0], b[158][1],b[158][2],b[158][3],b[158][4],b[158][5],b[158][6],b[158][7],b[158][8],b[158][9],b[158][10],b[158][11],b[158][12],b[158][13],b[158][14],b[158][15]}; 
{b[160][0], b[160][1],b[160][2],b[160][3],b[160][4],b[160][5],b[160][6],b[160][7],b[160][8],b[160][9],b[160][10],b[160][11],b[160][12],b[160][13],b[160][14],b[160][15]} <= {b[159][0], b[159][1],b[159][2],b[159][3],b[159][4],b[159][5],b[159][6],b[159][7],b[159][8],b[159][9],b[159][10],b[159][11],b[159][12],b[159][13],b[159][14],b[159][15]}; 
{b[161][0], b[161][1],b[161][2],b[161][3],b[161][4],b[161][5],b[161][6],b[161][7],b[161][8],b[161][9],b[161][10],b[161][11],b[161][12],b[161][13],b[161][14],b[161][15]} <= {b[160][0], b[160][1],b[160][2],b[160][3],b[160][4],b[160][5],b[160][6],b[160][7],b[160][8],b[160][9],b[160][10],b[160][11],b[160][12],b[160][13],b[160][14],b[160][15]}; 
{b[162][0], b[162][1],b[162][2],b[162][3],b[162][4],b[162][5],b[162][6],b[162][7],b[162][8],b[162][9],b[162][10],b[162][11],b[162][12],b[162][13],b[162][14],b[162][15]} <= {b[161][0], b[161][1],b[161][2],b[161][3],b[161][4],b[161][5],b[161][6],b[161][7],b[161][8],b[161][9],b[161][10],b[161][11],b[161][12],b[161][13],b[161][14],b[161][15]}; 
{b[163][0], b[163][1],b[163][2],b[163][3],b[163][4],b[163][5],b[163][6],b[163][7],b[163][8],b[163][9],b[163][10],b[163][11],b[163][12],b[163][13],b[163][14],b[163][15]} <= {b[162][0], b[162][1],b[162][2],b[162][3],b[162][4],b[162][5],b[162][6],b[162][7],b[162][8],b[162][9],b[162][10],b[162][11],b[162][12],b[162][13],b[162][14],b[162][15]}; 
{b[164][0], b[164][1],b[164][2],b[164][3],b[164][4],b[164][5],b[164][6],b[164][7],b[164][8],b[164][9],b[164][10],b[164][11],b[164][12],b[164][13],b[164][14],b[164][15]} <= {b[163][0], b[163][1],b[163][2],b[163][3],b[163][4],b[163][5],b[163][6],b[163][7],b[163][8],b[163][9],b[163][10],b[163][11],b[163][12],b[163][13],b[163][14],b[163][15]}; 
{b[165][0], b[165][1],b[165][2],b[165][3],b[165][4],b[165][5],b[165][6],b[165][7],b[165][8],b[165][9],b[165][10],b[165][11],b[165][12],b[165][13],b[165][14],b[165][15]} <= {b[164][0], b[164][1],b[164][2],b[164][3],b[164][4],b[164][5],b[164][6],b[164][7],b[164][8],b[164][9],b[164][10],b[164][11],b[164][12],b[164][13],b[164][14],b[164][15]}; 
{b[166][0], b[166][1],b[166][2],b[166][3],b[166][4],b[166][5],b[166][6],b[166][7],b[166][8],b[166][9],b[166][10],b[166][11],b[166][12],b[166][13],b[166][14],b[166][15]} <= {b[165][0], b[165][1],b[165][2],b[165][3],b[165][4],b[165][5],b[165][6],b[165][7],b[165][8],b[165][9],b[165][10],b[165][11],b[165][12],b[165][13],b[165][14],b[165][15]}; 
{b[167][0], b[167][1],b[167][2],b[167][3],b[167][4],b[167][5],b[167][6],b[167][7],b[167][8],b[167][9],b[167][10],b[167][11],b[167][12],b[167][13],b[167][14],b[167][15]} <= {b[166][0], b[166][1],b[166][2],b[166][3],b[166][4],b[166][5],b[166][6],b[166][7],b[166][8],b[166][9],b[166][10],b[166][11],b[166][12],b[166][13],b[166][14],b[166][15]}; 
{b[168][0], b[168][1],b[168][2],b[168][3],b[168][4],b[168][5],b[168][6],b[168][7],b[168][8],b[168][9],b[168][10],b[168][11],b[168][12],b[168][13],b[168][14],b[168][15]} <= {b[167][0], b[167][1],b[167][2],b[167][3],b[167][4],b[167][5],b[167][6],b[167][7],b[167][8],b[167][9],b[167][10],b[167][11],b[167][12],b[167][13],b[167][14],b[167][15]}; 
{b[169][0], b[169][1],b[169][2],b[169][3],b[169][4],b[169][5],b[169][6],b[169][7],b[169][8],b[169][9],b[169][10],b[169][11],b[169][12],b[169][13],b[169][14],b[169][15]} <= {b[168][0], b[168][1],b[168][2],b[168][3],b[168][4],b[168][5],b[168][6],b[168][7],b[168][8],b[168][9],b[168][10],b[168][11],b[168][12],b[168][13],b[168][14],b[168][15]}; 
{b[170][0], b[170][1],b[170][2],b[170][3],b[170][4],b[170][5],b[170][6],b[170][7],b[170][8],b[170][9],b[170][10],b[170][11],b[170][12],b[170][13],b[170][14],b[170][15]} <= {b[169][0], b[169][1],b[169][2],b[169][3],b[169][4],b[169][5],b[169][6],b[169][7],b[169][8],b[169][9],b[169][10],b[169][11],b[169][12],b[169][13],b[169][14],b[169][15]}; 
{b[171][0], b[171][1],b[171][2],b[171][3],b[171][4],b[171][5],b[171][6],b[171][7],b[171][8],b[171][9],b[171][10],b[171][11],b[171][12],b[171][13],b[171][14],b[171][15]} <= {b[170][0], b[170][1],b[170][2],b[170][3],b[170][4],b[170][5],b[170][6],b[170][7],b[170][8],b[170][9],b[170][10],b[170][11],b[170][12],b[170][13],b[170][14],b[170][15]}; 
{b[172][0], b[172][1],b[172][2],b[172][3],b[172][4],b[172][5],b[172][6],b[172][7],b[172][8],b[172][9],b[172][10],b[172][11],b[172][12],b[172][13],b[172][14],b[172][15]} <= {b[171][0], b[171][1],b[171][2],b[171][3],b[171][4],b[171][5],b[171][6],b[171][7],b[171][8],b[171][9],b[171][10],b[171][11],b[171][12],b[171][13],b[171][14],b[171][15]}; 
{b[173][0], b[173][1],b[173][2],b[173][3],b[173][4],b[173][5],b[173][6],b[173][7],b[173][8],b[173][9],b[173][10],b[173][11],b[173][12],b[173][13],b[173][14],b[173][15]} <= {b[172][0], b[172][1],b[172][2],b[172][3],b[172][4],b[172][5],b[172][6],b[172][7],b[172][8],b[172][9],b[172][10],b[172][11],b[172][12],b[172][13],b[172][14],b[172][15]}; 
{b[174][0], b[174][1],b[174][2],b[174][3],b[174][4],b[174][5],b[174][6],b[174][7],b[174][8],b[174][9],b[174][10],b[174][11],b[174][12],b[174][13],b[174][14],b[174][15]} <= {b[173][0], b[173][1],b[173][2],b[173][3],b[173][4],b[173][5],b[173][6],b[173][7],b[173][8],b[173][9],b[173][10],b[173][11],b[173][12],b[173][13],b[173][14],b[173][15]}; 
{b[175][0], b[175][1],b[175][2],b[175][3],b[175][4],b[175][5],b[175][6],b[175][7],b[175][8],b[175][9],b[175][10],b[175][11],b[175][12],b[175][13],b[175][14],b[175][15]} <= {b[174][0], b[174][1],b[174][2],b[174][3],b[174][4],b[174][5],b[174][6],b[174][7],b[174][8],b[174][9],b[174][10],b[174][11],b[174][12],b[174][13],b[174][14],b[174][15]}; 
{b[176][0], b[176][1],b[176][2],b[176][3],b[176][4],b[176][5],b[176][6],b[176][7],b[176][8],b[176][9],b[176][10],b[176][11],b[176][12],b[176][13],b[176][14],b[176][15]} <= {b[175][0], b[175][1],b[175][2],b[175][3],b[175][4],b[175][5],b[175][6],b[175][7],b[175][8],b[175][9],b[175][10],b[175][11],b[175][12],b[175][13],b[175][14],b[175][15]}; 
{b[177][0], b[177][1],b[177][2],b[177][3],b[177][4],b[177][5],b[177][6],b[177][7],b[177][8],b[177][9],b[177][10],b[177][11],b[177][12],b[177][13],b[177][14],b[177][15]} <= {b[176][0], b[176][1],b[176][2],b[176][3],b[176][4],b[176][5],b[176][6],b[176][7],b[176][8],b[176][9],b[176][10],b[176][11],b[176][12],b[176][13],b[176][14],b[176][15]}; 
{b[178][0], b[178][1],b[178][2],b[178][3],b[178][4],b[178][5],b[178][6],b[178][7],b[178][8],b[178][9],b[178][10],b[178][11],b[178][12],b[178][13],b[178][14],b[178][15]} <= {b[177][0], b[177][1],b[177][2],b[177][3],b[177][4],b[177][5],b[177][6],b[177][7],b[177][8],b[177][9],b[177][10],b[177][11],b[177][12],b[177][13],b[177][14],b[177][15]}; 
{b[179][0], b[179][1],b[179][2],b[179][3],b[179][4],b[179][5],b[179][6],b[179][7],b[179][8],b[179][9],b[179][10],b[179][11],b[179][12],b[179][13],b[179][14],b[179][15]} <= {b[178][0], b[178][1],b[178][2],b[178][3],b[178][4],b[178][5],b[178][6],b[178][7],b[178][8],b[178][9],b[178][10],b[178][11],b[178][12],b[178][13],b[178][14],b[178][15]}; 
{b[180][0], b[180][1],b[180][2],b[180][3],b[180][4],b[180][5],b[180][6],b[180][7],b[180][8],b[180][9],b[180][10],b[180][11],b[180][12],b[180][13],b[180][14],b[180][15]} <= {b[179][0], b[179][1],b[179][2],b[179][3],b[179][4],b[179][5],b[179][6],b[179][7],b[179][8],b[179][9],b[179][10],b[179][11],b[179][12],b[179][13],b[179][14],b[179][15]}; 
{b[181][0], b[181][1],b[181][2],b[181][3],b[181][4],b[181][5],b[181][6],b[181][7],b[181][8],b[181][9],b[181][10],b[181][11],b[181][12],b[181][13],b[181][14],b[181][15]} <= {b[180][0], b[180][1],b[180][2],b[180][3],b[180][4],b[180][5],b[180][6],b[180][7],b[180][8],b[180][9],b[180][10],b[180][11],b[180][12],b[180][13],b[180][14],b[180][15]}; 
{b[182][0], b[182][1],b[182][2],b[182][3],b[182][4],b[182][5],b[182][6],b[182][7],b[182][8],b[182][9],b[182][10],b[182][11],b[182][12],b[182][13],b[182][14],b[182][15]} <= {b[181][0], b[181][1],b[181][2],b[181][3],b[181][4],b[181][5],b[181][6],b[181][7],b[181][8],b[181][9],b[181][10],b[181][11],b[181][12],b[181][13],b[181][14],b[181][15]}; 
{b[183][0], b[183][1],b[183][2],b[183][3],b[183][4],b[183][5],b[183][6],b[183][7],b[183][8],b[183][9],b[183][10],b[183][11],b[183][12],b[183][13],b[183][14],b[183][15]} <= {b[182][0], b[182][1],b[182][2],b[182][3],b[182][4],b[182][5],b[182][6],b[182][7],b[182][8],b[182][9],b[182][10],b[182][11],b[182][12],b[182][13],b[182][14],b[182][15]}; 
{b[184][0], b[184][1],b[184][2],b[184][3],b[184][4],b[184][5],b[184][6],b[184][7],b[184][8],b[184][9],b[184][10],b[184][11],b[184][12],b[184][13],b[184][14],b[184][15]} <= {b[183][0], b[183][1],b[183][2],b[183][3],b[183][4],b[183][5],b[183][6],b[183][7],b[183][8],b[183][9],b[183][10],b[183][11],b[183][12],b[183][13],b[183][14],b[183][15]}; 
{b[185][0], b[185][1],b[185][2],b[185][3],b[185][4],b[185][5],b[185][6],b[185][7],b[185][8],b[185][9],b[185][10],b[185][11],b[185][12],b[185][13],b[185][14],b[185][15]} <= {b[184][0], b[184][1],b[184][2],b[184][3],b[184][4],b[184][5],b[184][6],b[184][7],b[184][8],b[184][9],b[184][10],b[184][11],b[184][12],b[184][13],b[184][14],b[184][15]}; 
{b[186][0], b[186][1],b[186][2],b[186][3],b[186][4],b[186][5],b[186][6],b[186][7],b[186][8],b[186][9],b[186][10],b[186][11],b[186][12],b[186][13],b[186][14],b[186][15]} <= {b[185][0], b[185][1],b[185][2],b[185][3],b[185][4],b[185][5],b[185][6],b[185][7],b[185][8],b[185][9],b[185][10],b[185][11],b[185][12],b[185][13],b[185][14],b[185][15]}; 
{b[187][0], b[187][1],b[187][2],b[187][3],b[187][4],b[187][5],b[187][6],b[187][7],b[187][8],b[187][9],b[187][10],b[187][11],b[187][12],b[187][13],b[187][14],b[187][15]} <= {b[186][0], b[186][1],b[186][2],b[186][3],b[186][4],b[186][5],b[186][6],b[186][7],b[186][8],b[186][9],b[186][10],b[186][11],b[186][12],b[186][13],b[186][14],b[186][15]}; 
{b[188][0], b[188][1],b[188][2],b[188][3],b[188][4],b[188][5],b[188][6],b[188][7],b[188][8],b[188][9],b[188][10],b[188][11],b[188][12],b[188][13],b[188][14],b[188][15]} <= {b[187][0], b[187][1],b[187][2],b[187][3],b[187][4],b[187][5],b[187][6],b[187][7],b[187][8],b[187][9],b[187][10],b[187][11],b[187][12],b[187][13],b[187][14],b[187][15]}; 
{b[189][0], b[189][1],b[189][2],b[189][3],b[189][4],b[189][5],b[189][6],b[189][7],b[189][8],b[189][9],b[189][10],b[189][11],b[189][12],b[189][13],b[189][14],b[189][15]} <= {b[188][0], b[188][1],b[188][2],b[188][3],b[188][4],b[188][5],b[188][6],b[188][7],b[188][8],b[188][9],b[188][10],b[188][11],b[188][12],b[188][13],b[188][14],b[188][15]}; 
{b[190][0], b[190][1],b[190][2],b[190][3],b[190][4],b[190][5],b[190][6],b[190][7],b[190][8],b[190][9],b[190][10],b[190][11],b[190][12],b[190][13],b[190][14],b[190][15]} <= {b[189][0], b[189][1],b[189][2],b[189][3],b[189][4],b[189][5],b[189][6],b[189][7],b[189][8],b[189][9],b[189][10],b[189][11],b[189][12],b[189][13],b[189][14],b[189][15]}; 
{b[191][0], b[191][1],b[191][2],b[191][3],b[191][4],b[191][5],b[191][6],b[191][7],b[191][8],b[191][9],b[191][10],b[191][11],b[191][12],b[191][13],b[191][14],b[191][15]} <= {b[190][0], b[190][1],b[190][2],b[190][3],b[190][4],b[190][5],b[190][6],b[190][7],b[190][8],b[190][9],b[190][10],b[190][11],b[190][12],b[190][13],b[190][14],b[190][15]}; 
{b[192][0], b[192][1],b[192][2],b[192][3],b[192][4],b[192][5],b[192][6],b[192][7],b[192][8],b[192][9],b[192][10],b[192][11],b[192][12],b[192][13],b[192][14],b[192][15]} <= {b[191][0], b[191][1],b[191][2],b[191][3],b[191][4],b[191][5],b[191][6],b[191][7],b[191][8],b[191][9],b[191][10],b[191][11],b[191][12],b[191][13],b[191][14],b[191][15]}; 
{b[193][0], b[193][1],b[193][2],b[193][3],b[193][4],b[193][5],b[193][6],b[193][7],b[193][8],b[193][9],b[193][10],b[193][11],b[193][12],b[193][13],b[193][14],b[193][15]} <= {b[192][0], b[192][1],b[192][2],b[192][3],b[192][4],b[192][5],b[192][6],b[192][7],b[192][8],b[192][9],b[192][10],b[192][11],b[192][12],b[192][13],b[192][14],b[192][15]}; 
{b[194][0], b[194][1],b[194][2],b[194][3],b[194][4],b[194][5],b[194][6],b[194][7],b[194][8],b[194][9],b[194][10],b[194][11],b[194][12],b[194][13],b[194][14],b[194][15]} <= {b[193][0], b[193][1],b[193][2],b[193][3],b[193][4],b[193][5],b[193][6],b[193][7],b[193][8],b[193][9],b[193][10],b[193][11],b[193][12],b[193][13],b[193][14],b[193][15]}; 
{b[195][0], b[195][1],b[195][2],b[195][3],b[195][4],b[195][5],b[195][6],b[195][7],b[195][8],b[195][9],b[195][10],b[195][11],b[195][12],b[195][13],b[195][14],b[195][15]} <= {b[194][0], b[194][1],b[194][2],b[194][3],b[194][4],b[194][5],b[194][6],b[194][7],b[194][8],b[194][9],b[194][10],b[194][11],b[194][12],b[194][13],b[194][14],b[194][15]}; 
{b[196][0], b[196][1],b[196][2],b[196][3],b[196][4],b[196][5],b[196][6],b[196][7],b[196][8],b[196][9],b[196][10],b[196][11],b[196][12],b[196][13],b[196][14],b[196][15]} <= {b[195][0], b[195][1],b[195][2],b[195][3],b[195][4],b[195][5],b[195][6],b[195][7],b[195][8],b[195][9],b[195][10],b[195][11],b[195][12],b[195][13],b[195][14],b[195][15]}; 
{b[197][0], b[197][1],b[197][2],b[197][3],b[197][4],b[197][5],b[197][6],b[197][7],b[197][8],b[197][9],b[197][10],b[197][11],b[197][12],b[197][13],b[197][14],b[197][15]} <= {b[196][0], b[196][1],b[196][2],b[196][3],b[196][4],b[196][5],b[196][6],b[196][7],b[196][8],b[196][9],b[196][10],b[196][11],b[196][12],b[196][13],b[196][14],b[196][15]}; 
{b[198][0], b[198][1],b[198][2],b[198][3],b[198][4],b[198][5],b[198][6],b[198][7],b[198][8],b[198][9],b[198][10],b[198][11],b[198][12],b[198][13],b[198][14],b[198][15]} <= {b[197][0], b[197][1],b[197][2],b[197][3],b[197][4],b[197][5],b[197][6],b[197][7],b[197][8],b[197][9],b[197][10],b[197][11],b[197][12],b[197][13],b[197][14],b[197][15]}; 
{b[199][0], b[199][1],b[199][2],b[199][3],b[199][4],b[199][5],b[199][6],b[199][7],b[199][8],b[199][9],b[199][10],b[199][11],b[199][12],b[199][13],b[199][14],b[199][15]} <= {b[198][0], b[198][1],b[198][2],b[198][3],b[198][4],b[198][5],b[198][6],b[198][7],b[198][8],b[198][9],b[198][10],b[198][11],b[198][12],b[198][13],b[198][14],b[198][15]};
		i = 199;
		end
		else
		i = i + 1;
	 end
	 
endmodule
